library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY Reg_n IS
GENERIC(N: INTEGER :=9);
PORT(
	CLK, RST_n: IN STD_LOGIC;
	DIN: IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	DOUT: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END ENTITY; 

ARCHITECTURE beh OF Reg_n IS 
	
BEGIN
	PROCESS(CLK)
	BEGIN
		IF CLK'EVENT AND CLK = '1' THEN
			IF RST_n = '0' THEN
				DOUT <= (OTHERS => '0');
			ELSE
				DOUT <= DIN;
			END IF;
		END IF;
	END PROCESS;
END beh;